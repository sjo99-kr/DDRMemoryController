`timescale 1ns / 1ps

//------------------------------------------------------------------------------
//      RankSched
//
//      Role:
//          Rank-level request scheduler for DDR memory system.
//
//      Responsibilities:
//          - Buffers read/write requests from MC frontend.
//          - Applies FR-FCFS policy with open-page awareness.
//          - Manages refresh scheduling (tREFI).
//          - Selects next request to issue to RankFSM.
//          - Tracks open rows and request aging.
//
//      Scheduling Policy:
//          - FR-FCFS (First-Ready, First-Come-First-Serve)
//          - Priority order:
//              1) Requests beyond aging threshold
//              2) Row-hit with short tCCD
//              3) Row-hit with long tCCD
//              4) Oldest request (aging-based)
//
//      Scope & Notes:
//          - Operates at rank granularity.
//          - No command-level timing (handled by RankFSM).
//          - One request issued at a time to RankFSM.
//
//      Author  : Seongwon Jo
//      Created : 2026.02
//------------------------------------------------------------------------------
import MemoryController_Definitions::*;

module RankSched (
    // Common
    input logic clk, rst,

    input [32-1:0] RankReqMemAddr,                                             
    input logic [MEM_IDWIDTH-1:0] RankReqId,                                 
    input logic [MEM_USERWIDTH-1:0] RankReqUser,                            
    input logic RankReqType, 
    input logic RankReqValid,                              
                     
    output logic RankReadReqReady,                    // Valid When RD Req. Que. is not full & RD MEM Buffer is available
    output logic RankWriteReqReady,                   // Valid When WR Req. Que. is not full & WR MEM Buffer is available

                                                          //   Input from Channel Scheduler    //
    input logic chSchedCMDOnlyValid,                  //  (Input from Channel Scheduler)   //
    input logic chSchedCMDDQValid,                    //  (Input from Channel Scheduler)   //
    input wire chSchedTransReady,
    output logic chSchedAvailableCMD,                 //       (Output to RankFSM)         //
    output logic chSchedAvailableCMDDQ,                //       (Output to RankFSM)         //

    input logic WriteMode,                            

    output logic chSchedRdReady,      
    output logic chSchedWrReady,

    input logic fsmChSchedAck,                        //      (Input from RankFSM)         //    
    input logic [NUM_BANKFSM-1:0] fsmWait,                              //      (Input fron RankFSM)         //
                                                          //  Valid when RankFSM is WAITING for DRAM TIMING CONSTRAINTS.    
    output logic chSchedACK,                          //       (Output to RankFSM)         //
    output logic chSchedIdle,                         //       (Output to RankFSM)         //
        
    output logic [$clog2(READCMDQUEUEDEPTH)-1:0] chSchedReadReqCnt,
    output logic [$clog2(WRITECMDQUEUEDEPTH)-1:0] chSchedWriteReqCnt,

    input logic rdBufAvailable,                       //    (Input from MEM Buffer)      //
    input logic wrBufAvailable,                       //    (Input from MEM Buffer)      //
    output logic fsmWrBufValid,                       //        (Ouput to RankFSM)       //
    output logic fsmRdBufValid,                       //        (Ouput to RankFSM)       //

    output logic [MEM_IDWIDTH-1:0] readBufReqId, 
    output logic [MEM_USERWIDTH-1:0] readBufReqUser,
    output logic readBufReqACK,
    output logic [MEM_IDWIDTH-1:0] writeBufReqId,
    output logic [MEM_USERWIDTH-1:0] writeBufReqUser,
    output logic writeBufReqACK,

    input logic [NUM_BANKFSM-1:0] fsmIdle,                              // Valid when RankFSM is Idle State, Ready for receiving NEW REQUEST.
    input logic fsmRefreshAck,                        // Valid when RankFSM finished Refresh phase.
    output logic refresh,                             // Valid when the timing for tREFI is set.

    input logic [MEM_IDWIDTH-1:0] fsmBufWrReqId, fsmBufRdReqId,
    input logic [MEM_USERWIDTH-1:0] fsmBufWrReqUser, fsmBufRdReqUser, 
    input logic fsmBufWrReqIssued,                 
    input logic fsmBufRdReqIssued,

    output logic [NUM_BANKFSM-1:0] fsmIssue,                            // Valid when Request Scheduler sends Request to RankFSM.
    output [44-1:0] fsmIssuedReq,                       // Request for RankFSM when RankFSM is Idle.
    output logic issuable
    );

    localparam int CMDQUEUEDEPTH = (READCMDQUEUEDEPTH > WRITECMDQUEUEDEPTH) ? READCMDQUEUEDEPTH : WRITECMDQUEUEDEPTH;

    //------------------------ Interface signals Setup ----------------------//
    //                RankSched/FSM <-> ChannelSched/Arbiter                 //
    assign chSchedRdReady =  !fsmIdle && !fsmWait; // 이거 다시 시그널 설정하기!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
    assign chSchedWrReady =  !fsmIdle && !fsmWait; // 이거 다시 시그널 설정하기!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
    assign chSchedIdle = fsmWait;
    assign chSchedACK = fsmChSchedAck;                  

    assign chSchedAvailableCMD = chSchedCMDOnlyValid;
    assign chSchedAvailableCMDDQ = chSchedCMDDQValid;

    //                  MEMBuffer-side <-> RankSched/FSM                   //
    assign readBufReqId = fsmBufRdReqId;
    assign readBufReqUser = fsmBufRdReqUser;

    assign writeBufReqId = fsmBufWrReqId;
    assign writeBufReqUser = fsmBufWrReqUser;

    assign writeBufReqACK = fsmBufWrReqIssued;
    assign readBufReqACK = fsmBufRdReqIssued;

    assign fsmRdBufValid = rdBufAvailable;
    assign fsmWrBufValid = wrBufAvailable;
    //////////////////////////////////////////////////////////////////////////

    //------------------------ Struct Definition ---------------------------//
    typedef struct packed{
        logic[32-1:0] mem_addr;  // [47:16]
        logic req_type; // [15]
        logic [MEM_IDWIDTH-1:0] req_id; // [14]
        logic [MEM_USERWIDTH-1:0] req_user;  // [13:10]
        logic [AGINGWIDTH-1:0] cnt; // [9:0]
    } ReqQueEntry; // 48

    typedef struct packed {
        logic valid;
        logic [RWIDTH-1:0] RowAddr;
    }OpenRowEntry;
    //////////////////////////////////////////////////////////////////////////

    //      Memory Request Queue for Read Request and Write Request         //
    ReqQueEntry [0: READCMDQUEUEDEPTH - 1] ReadRequestQueue;
    ReqQueEntry [0: WRITECMDQUEUEDEPTH - 1] WriteRequestQueue;
    logic [$clog2(READCMDQUEUEDEPTH) - 1 : 0] ReadPushPtr, ReadPopPtr;
    logic [$clog2(WRITECMDQUEUEDEPTH) - 1 : 0] WritePushPtr, WritePopPtr;
    logic [READCMDQUEUEDEPTH - 1:0] ReadReqQueFree;
    logic [WRITECMDQUEUEDEPTH - 1:0] WriteReqQueFree;
    logic ReadReqQueFull, ReadReqQueEmpty; 
    logic WriteReqQueFull, WriteReqQueEmpty;

    //            OpenPagePolicy management  (OpenPagePolicy List)         //
    OpenRowEntry OpenRowList [OPENPAGELISTDEPTH - 1 : 0 ];              // OpenRowDepth -> Num. of BankGroup * Num. of Bank., One bank has one Row (Page).
    logic checkThreshold;                                          // Threshold for blocking starvation in Request Queue. (request aging)
    logic [$clog2(CMDQUEUEDEPTH) - 1 : 0] MaxValue;                  // MaxValue for Oldes Entry in Request Queue.
    
    logic [1:0] PageHitT;                                          // PageHit indicates a row-hit condition within a bank.
                                                                   // In a row-hit case, READ or WRITE commands can be issued
                                                                   // without an ACT command.
                                                                   //
                                                                   // When consecutive column commands (READ/WRITE) are issued:
                                                                   // - If the commands target banks within the same bank group,
                                                                   //    tCCD_S (short) timing constraint applies.
                                                                   // - If the commands target banks in different bank groups,
                                                                   //    tCCD_L (long) timing constraint applies.

    logic PageMissT, PageEmptyT;                                   // PageMiss -> Need to Precharge on current Row(Page), and ACT the target Row.
                                                                   // PageEmpty -> Need to ACT the target Row without Precharge
    logic NextPageHitS, NextPageHitL;       
    logic [$clog2(CMDQUEUEDEPTH) -1 :0] PageHitIndexS, PageHitIndexL;

    // Refresh management
    logic [$clog2(tREFI)-1:0] refresh_cnt;                         // Refresh Interval Count
    logic refreshing;                                              // Refresh flag.
                                                                   // Normally, refresh is issued at the rank level.

    // AutoPrecharge Commnad
    logic checkAutoPrecharge;

    //------------------------------------------------------------------------------
    //  Refresh Scheduler
    //
    //  - Tracks refresh interval (tREFI).
    //  - Issues rank-level refresh request when interval expires.
    //  - Refresh is only triggered when RankFSM is idle.
    //
    //------------------------------------------------------------------------------
    always_ff@(posedge clk or negedge rst)begin
        if(!rst) begin
            refresh_cnt <= 0;
            refreshing <= 0;
        end else begin
            if(refreshing == 0) begin
                refresh_cnt <= refresh_cnt + 1;
                if(refresh_cnt == (tREFI - 1)) begin        // tREFI : Refresh Interval Cycles.
                    refreshing <= 1;                        // Refresh Flag Setup.
                    refresh_cnt <= 0;
                end
            end else begin
                if(fsmRefreshAck) begin                     // ACK from RankFSM for Refreshing done.
                    refreshing <= 0; 
                end
            end
        end
    end
    assign refresh = refreshing;            // Refresh send when RankFSM is IDLE.  
                                                            // (TODO) : Refresh needs to be availble whenever the flag is set on.
    //////////////////////////////////////////////////////////////////////////


    //------------------------------------------------------------------------------
    //  Request Count Export
    //
    //  - Counts outstanding read/write requests in queues.
    //  - Used by ChannelScheduler for arbitration decisions.
    //
    //------------------------------------------------------------------------------
    always_comb begin
        chSchedReadReqCnt = 0;
        chSchedWriteReqCnt = 0;
        for(int i = 0; i < READCMDQUEUEDEPTH; i++) begin
            if(!ReadReqQueFree[i]) begin
                chSchedReadReqCnt = chSchedReadReqCnt + 1;
            end
        end
        for (int i = 0; i < WRITECMDQUEUEDEPTH; i++) begin
            if(!WriteReqQueFree[i]) begin
                chSchedWriteReqCnt = chSchedWriteReqCnt + 1;
            end
        end
    end
    //////////////////////////////////////////////////////////////////////////

    //------------------ Memory Request Queue Setup ------------------------//
    //               Set up Push Pointer based on LSB priority              //
    PriorityEncoder_LSB push_ptr(     
        .vector(ReadReqQueFree),
        .index(ReadPushPtr)
    );

    PriorityEncoder_LSB  write_push_ptr( 
        .vector(WriteReqQueFree),
        .index(WritePushPtr)
    );

    //------------------------------------------------------------------------------
    //  Request Queue Management
    //
    //  - Pushes incoming requests from MC frontend.
    //  - Pops selected request when RankFSM is idle.
    //  - Maintains free-slot bitmap and push/pop pointers.
    //  - Includes structural hazard assertions.
    //
    //------------------------------------------------------------------------------
    always_ff@(posedge clk or negedge rst) begin
        if(!rst)begin
             // Free Queue Setup, 1 for Free slot, 0 for Allocated slot
            ReadReqQueFree <= '1;             
            WriteReqQueFree <= '1;
            //  Read/Write Request Queue Initialization (without count)
            for(int i = 0; i < READCMDQUEUEDEPTH; i++) begin
                ReadRequestQueue[i][47:16] <= 0;
                ReadRequestQueue[i][15] <= 0;
                ReadRequestQueue[i][14] <= 0;
                ReadRequestQueue[i][13:10] <= 0;
            end
            for(int i = 0; i < WRITECMDQUEUEDEPTH; i++) begin
                WriteRequestQueue[i][47:16] <= 0;
                WriteRequestQueue[i][15] <= 0;
                WriteRequestQueue[i][14] <= 0;
                WriteRequestQueue[i][13:10] <= 0;
            end
        end else begin
            //          Push Phase: Pushing Req. from MC FrontEnd           //
            if(RankReqValid && !ReadReqQueFull && (RankReqType == 0)) begin
                // For Read Request Case
                ReadRequestQueue[ReadPushPtr][47:16] <= RankReqMemAddr;
                ReadRequestQueue[ReadPushPtr][15] <= RankReqType;
                ReadRequestQueue[ReadPushPtr][14] <= RankReqId;
                ReadRequestQueue[ReadPushPtr][13:10] <= RankReqUser;
                ReadReqQueFree[ReadPushPtr] <= 0;
            end
            if(RankReqValid && !WriteReqQueFull && (RankReqType == 1)) begin
                // For Write Request Case
                WriteRequestQueue[WritePushPtr][47:16] <= RankReqMemAddr;
                WriteRequestQueue[WritePushPtr][15] <= RankReqType;
                WriteRequestQueue[WritePushPtr][14] <= RankReqId;
                WriteRequestQueue[WritePushPtr][13:10] <= RankReqUser;
                WriteReqQueFree[WritePushPtr] <= '0;
            end
            //     POP Phase: Poping Req. Request Que. and send to RankFSM   //
            if(fsmIdle[{ReadRequestQueue[ReadPopPtr][40:39], ReadRequestQueue[ReadPopPtr][38:37]}]
                 && !ReadReqQueFree[ReadPopPtr] && !WriteMode && !refreshing && !chSchedTransReady) begin 
                // For Read Request Case (Initialization for Request Queue)
                ReadRequestQueue[ReadPopPtr][47:16] <= 0; 
                ReadRequestQueue[ReadPopPtr][15] <= 0;
                ReadRequestQueue[ReadPopPtr][14] <= 0;
                ReadRequestQueue[ReadPopPtr][13:10] <= 0;
                ReadReqQueFree[ReadPopPtr] <= '1;
            end 
            if(fsmIdle[{WriteRequestQueue[WritePopPtr][40:39], WriteRequestQueue[WritePopPtr][38:37]}]
                && !WriteReqQueFree[WritePopPtr] && WriteMode && !refreshing && !chSchedTransReady) begin
                // For Write Request Case (Initialization for Request Queue)
                WriteRequestQueue[WritePopPtr][47:16] <= 0; 
                WriteRequestQueue[WritePopPtr][15] <= 0;
                WriteRequestQueue[WritePopPtr][14] <= 0;
                WriteRequestQueue[WritePopPtr][13:10] <= 0;
                WriteReqQueFree[WritePopPtr] <= '1;
            end
        end
    end

    assign ReadReqQueFull = !(|ReadReqQueFree);
    assign ReadReqQueEmpty = (&ReadReqQueFree);
    assign WriteReqQueFull = !(|WriteReqQueFree);
    assign WriteReqQueEmpty = (&WriteReqQueFree);

    assign RankReadReqReady =  !ReadReqQueFull && rdBufAvailable;
    assign RankWriteReqReady = !WriteReqQueFull && wrBufAvailable;


    //------------------------------------------------------------------------------
    //  Request Aging Tracker
    //
    //  - Increments per-request age counters.
    //  - Resets age when request is issued to RankFSM.
    //  - Enables starvation prevention via threshold logic.
    //
    //------------------------------------------------------------------------------
        always_ff@(posedge clk or negedge rst)begin
        // Request Count Setup for aging
        if(!rst) begin
            for(int i = 0; i < READCMDQUEUEDEPTH; i++) begin
                ReadRequestQueue[i][9:0] <= 0;
            end
            for (int i = 0; i< WRITECMDQUEUEDEPTH; i++) begin
                WriteRequestQueue[i][9:0] <= 0;
            end
        end else begin
            for(int i = 0; i < READCMDQUEUEDEPTH; i++)begin
                if(!ReadReqQueFree[i]) begin
                    ReadRequestQueue[i][9:0] <= ReadRequestQueue[i][9:0] + 1;
                end
            end
            for(int i = 0; i < WRITECMDQUEUEDEPTH; i++) begin
                if(!WriteReqQueFree[i]) begin
                    WriteRequestQueue[i][9:0] <= WriteRequestQueue[i][9:0] + 1; 
                end
            end
            if(fsmIdle && !ReadReqQueFree[ReadPopPtr] && !WriteMode && !refreshing) begin // Condition for Sending Req. to RankFSM
                ReadRequestQueue[ReadPopPtr][9:0] <= 0;
            end
            if(fsmIdle && !WriteReqQueFree[WritePopPtr] && WriteMode && !refreshing) begin // Condition for Sending Req. to RankFSM
                WriteRequestQueue[WritePopPtr][9:0] <= 0;
            end

        end
    end
    //////////////////////////////////////////////////////////////////////////
    

    //------------------------------------------------------------------------------
    //  RankFSM Issue Logic & Open-Page Update
    //
    //  - Issues selected request to RankFSM.
    //  - Updates OpenRowList on ACT / Auto-Precharge.
    //  - Clears open-page state on refresh completion.
    //
    //------------------------------------------------------------------------------
    always_ff@(posedge clk or negedge rst) begin
        if(!rst) begin
            fsmIssuedReq <= '0;                 //  Request to RankFSM
            for(int j = 0; j < NUM_BANKFSM; j++) begin
                fsmIssue[j] <= 0;               //  Valid when issuing REQUEST to RankFSM
            end
            for(int i = 0; i < OPENPAGELISTDEPTH; i++)begin
                OpenRowList[i] <= '0;           // Initialization of OpenRowList
            end  
        end else begin 
            if(fsmRefreshAck) begin             // Initialization of OpenRowList, when Refresh ACK comes on.
                                                // - Refresh is executed after precharging all pages, so we need to initialize OpenRowList.
                for(int i = 0; i < OPENPAGELISTDEPTH; i++) begin
                    OpenRowList[i] <= '0;
                end
            end
            if (!chSchedTransReady && !refreshing) begin                           // Sending Request to RankFSM based on the Condition.
                if(fsmIdle[{ReadRequestQueue[ReadPopPtr][40:39], ReadRequestQueue[ReadPopPtr][38:37]}] &&
                !WriteMode && !ReadReqQueFree[ReadPopPtr]) begin 
                    fsmIssuedReq[43:12] <= ReadRequestQueue[ReadPopPtr][43:12];
                    fsmIssuedReq[5] <= ReadRequestQueue[ReadPopPtr][5];
                    {fsmIssuedReq[11:9], fsmIssuedReq[8], fsmIssuedReq[7]} <= {PageHitT, PageMissT, PageEmptyT};
                    fsmIssuedReq[4] <= ReadRequestQueue[ReadPopPtr][4];
                    fsmIssuedReq[3:0] <= ReadRequestQueue[ReadPopPtr][3:0];
                    fsmIssue[{ReadRequestQueue[ReadPopPtr][40:39], ReadRequestQueue[ReadPopPtr][38:37]}] <= 1;
                    $display("[CH-%d RK-%D SCHED] CLK: %d | READ REQUEST SEND", FSM_CHANNEL, FSM_RANK, $time);

                    //           For AutoPrecharge Instruction, we invalidate AutoPrecharge Page in OpenPageList.            //
                    if(!checkAutoPrecharge) begin
                        //      If the Request is not for AutoPrecharge, then we just allocate that request in OpenPageList     //
                        OpenRowList[{ReadRequestQueue[ReadPopPtr][40:39], ReadRequestQueue[ReadPopPtr][38:37]}][15] <= 1;
                        OpenRowList[{ReadRequestQueue[ReadPopPtr][40:39], ReadRequestQueue[ReadPopPtr][38:37]}][14:0] <=
                            ReadRequestQueue[ReadPopPtr][36:22];
                        fsmIssuedReq[6] <= 0;
                    end else begin
                        OpenRowList[{ReadRequestQueue[ReadPopPtr][40:39], ReadRequestQueue[ReadPopPtr][38:37]}][15] <= 0;
                        fsmIssuedReq[6] <= 1;
                    end
                end else if(fsmIdle[{WriteRequestQueue[WritePopPtr][40:39], WriteRequestQueue[WritePopPtr][38:37]}] && 
                    WriteMode && !WriteReqQueFree[WritePopPtr]) begin
                    // Write Request Serving
                    fsmIssuedReq.mem_addr <= WriteRequestQueue[WritePopPtr][43:12];
                    fsmIssuedReq.req_type <= WriteRequestQueue[WritePopPtr][5];
                    {fsmIssuedReq[11:9], fsmIssuedReq[8], fsmIssuedReq[7]} <= {PageHitT, PageMissT, PageEmptyT};
                    fsmIssuedReq.req_user <= WriteRequestQueue[WritePopPtr][4];
                    fsmIssuedReq.req_id <= WriteRequestQueue[WritePopPtr][3:0];
                    fsmIssue[{WriteRequestQueue[WritePopPtr][40:39], WriteRequestQueue[WritePopPtr][38:37]}] <= 1;
                    $display("[CH-%d RK-%D SCHED] CLK: %d | WRITE REQUEST SEND", FSM_CHANNEL, FSM_RANK, $time);
                    //           For AutoPrecharge Instruction, we invalidate AutoPrecharge Page in OpenPageList.            //
                    if(!checkAutoPrecharge) begin
                        OpenRowList[{ReadRequestQueue[WritePopPtr][40:39], ReadRequestQueue[WritePopPtr][38:37]}][15] <= 1;
                        OpenRowList[{ReadRequestQueue[WritePopPtr][40:39], ReadRequestQueue[WritePopPtr][38:37]}][14:0] <=
                            ReadRequestQueue[WritePopPtr][36:22];
                        fsmIssuedReq[6] <= 0;
                    end else begin
                        OpenRowList[{ReadRequestQueue[WritePopPtr][40:39], ReadRequestQueue[WritePopPtr][38:37]}][15] <= 0;
                        fsmIssuedReq[6] <= 1;
                    end
                end else begin
                    for(int i = 0; i < NUM_BANKFSM; i++) begin
                        fsmIssue[i] <= 0;
                    end
                end
            end else begin
                for(int i = 0; i < NUM_BANKFSM; i++) begin
                    fsmIssue[i] <= 0;
                end
            end
        end
    end
    //////////////////////////////////////////////////////////////////////////

    logic issuableCheck, readIssuable, writeIssuable;
    assign issuableCheck =  (!refreshing && !chSchedTransReady);
    assign readIssuable = fsmIdle[{ReadRequestQueue[ReadPopPtr][40:39], ReadRequestQueue[ReadPopPtr][38:37]}] &&
                !WriteMode && !ReadReqQueFree[ReadPopPtr];

    assign writeIssuable = fsmIdle[{WriteRequestQueue[WritePopPtr][40:39], WriteRequestQueue[WritePopPtr][38:37]}] && 
                    WriteMode && !WriteReqQueFree[WritePopPtr];
                

    assign issuable = (WriteMode) ? writeIssuable : readIssuable;

    //------------------------------------------------------------------------------
    //  Open-Page Policy Helpers
    //
    //  - Detect row-hit candidates for short / long tCCD cases.
    //  - Separates same-bankgroup vs cross-bankgroup conditions.
    //  - Used by FR-FCFS candidate selection logic.
    //
    //------------------------------------------------------------------------------

    function automatic logic ReadOpenPagePolicyShort;
        input integer i;  // or input int i;
        begin
            if (
                ReadRequestQueue[i][36:22] ==
                OpenRowList[{ReadRequestQueue[i][40:39],
                             ReadRequestQueue[i][38:37]}][14:0]
                &&
                OpenRowList[{ReadRequestQueue[i][40:39],
                             ReadRequestQueue[i][38:37]}][15]
                &&
                !ReadReqQueFree[i]
                &&
                fsmIssuedReq[40:39] ==
                ReadRequestQueue[i][40:39]
            ) begin
                ReadOpenPagePolicyShort = 1'b1;
            end else begin
                ReadOpenPagePolicyShort = 1'b0;
            end
        end
    endfunction

        //////////////////////        Condition for Open for Short tCCD               /////////////////////
        // 1) Row Hit : Row of the target Request in Request Queue is SAME with the row in OpenPageList. //
        // 2) Request Valid : Request in Request Queue is valid for sending to RankFSM                   //
        // 3) Diff BG with Prior Req. : BankGroup (BG) of target Req is NOT SAME with BG with Prior Req. //
        ///////////////////////////////////////////////////////////////////////////////////////////////////
    function automatic logic ReadOpenPagePolicyLong;
        input integer i;
        begin
            if (
                (ReadRequestQueue[i][36:22] ==
                 OpenRowList[{ReadRequestQueue[i][40:39],
                              ReadRequestQueue[i][38:37]}][14:0])
                &&
                OpenRowList[{ReadRequestQueue[i][40:39],
                             ReadRequestQueue[i][38:37]}][15]
                &&
                !ReadReqQueFree[i]
                &&
                fsmIssuedReq[40:39] !=
                ReadRequestQueue[i][40:39]
            ) begin
                ReadOpenPagePolicyLong = 1'b1;
            end else begin
                ReadOpenPagePolicyLong = 1'b0;
            end
        end
    endfunction

//                    Write Request OpenPage Scheduling                 //
    function automatic logic WriteOpenPagePolicyShort;
        input integer i;
        begin
            if (
                WriteRequestQueue[i][36:22] ==
                OpenRowList[{WriteRequestQueue[i][40:39],
                             WriteRequestQueue[i][38:37]}][14:0]
                &&
                OpenRowList[{WriteRequestQueue[i][40:39],
                             WriteRequestQueue[i][38:37]}][15]
                &&
                !WriteReqQueFree[i]
                &&
                fsmIssuedReq[40:39] ==
                WriteRequestQueue[i][40:39]
            ) begin
                WriteOpenPagePolicyShort = 1'b1;
            end else begin
                WriteOpenPagePolicyShort = 1'b0;
            end
        end
    endfunction
    
    function automatic logic WriteOpenPagePolicyLong;
        input integer i;
        begin
            if (
                (WriteRequestQueue[i][36:22] ==
                 OpenRowList[{WriteRequestQueue[i][40:39],
                              WriteRequestQueue[i][38:37]}][14:0])
                &&
                OpenRowList[{WriteRequestQueue[i][40:39],
                             WriteRequestQueue[i][38:37]}][15]
                &&
                !WriteReqQueFree[i]
                &&
                (fsmIssuedReq[40:39] !=
                 WriteRequestQueue[i][40:39])
            ) begin
                WriteOpenPagePolicyLong = 1'b1;
            end else begin
                WriteOpenPagePolicyLong = 1'b0;
            end
        end
    endfunction
    //////////////////////////////////////////////////////////////////////////

    //------------------------------------------------------------------------------
    //  FR-FCFS Candidate Detection
    //
    //  - Identifies:
    //      * Short tCCD row-hits
    //      * Long tCCD row-hits
    //      * Oldest request (aging-based)
    //  - Separates read and write scheduling paths.
    //
    //------------------------------------------------------------------------------
    //        Candidate 1: Row Hit with Short-tCCD    PRIORITY: 2           //
    always_comb begin  
        NextPageHitS = 0;
        PageHitIndexS = '0;
        if(!WriteMode) begin
            // read request serving
            for(int i = READCMDQUEUEDEPTH-1; i>=0; i--)begin 
                if(ReadOpenPagePolicyShort(i) &&
                !fsmWait[{ReadRequestQueue[i][40:39], ReadRequestQueue[i][38:37]}] &&
                 fsmIdle[{ReadRequestQueue[i][40:39], ReadRequestQueue[i][38:37]}]
                 )begin
                    NextPageHitS = 1;
                    PageHitIndexS = i;
                end
            end
        end else begin
            // write request serving
            for(int i = WRITECMDQUEUEDEPTH-1; i>=0; i--) begin
                if(WriteOpenPagePolicyShort(i) &&
                !fsmWait[{WriteRequestQueue[i][40:39], WriteRequestQueue[i][38:37]}] &&
                 fsmIdle[{WriteRequestQueue[i][40:39], WriteRequestQueue[i][38:37]}]) 
                 begin
                    NextPageHitS = 1;
                    PageHitIndexS = i;
                end
            end
        end
    end
    //        Candidate 2: Row Hit with Long-tCCD     PRIORITY: 3         //
    always_comb begin 
        NextPageHitL = 0;
        PageHitIndexL = 0;
        if(!WriteMode) begin
            for(int i = READCMDQUEUEDEPTH-1; i>= 0; i--) begin
                if(ReadOpenPagePolicyLong(i) && 
                !fsmWait[{ReadRequestQueue[i][40:39], ReadRequestQueue[i][38:37]}] &&
                 fsmIdle[{ReadRequestQueue[i][40:39], ReadRequestQueue[i][38:37]}])
                 begin
                    NextPageHitL = 1;
                    PageHitIndexL = i[$clog2(READCMDQUEUEDEPTH)-1:0];
                end
            end
        end else begin
            for(int i = WRITECMDQUEUEDEPTH-1; i>=0; i--) begin
                if(WriteOpenPagePolicyLong(i) && 
                !fsmWait[{WriteRequestQueue[i][40:39], WriteRequestQueue[i][38:37]}] &&
                 fsmIdle[{WriteRequestQueue[i][40:39], WriteRequestQueue[i][38:37]}]
                 )begin
                    NextPageHitL = 1;
                    PageHitIndexL = i[$clog2(WRITECMDQUEUEDEPTH)-1:0];;
                end
            end
        end
    end

    //   Candidate 3: Under NO PAGEHIT, Oldest Request   PRIORITY: 4 (1)  //
    always_comb begin 
        MaxValue = 0;
        if(!WriteMode)begin
            // Read Request serving
            for(int i =0; i < READCMDQUEUEDEPTH; i++) begin
                if(!ReadReqQueFree[i] && (ReadRequestQueue[i][9:0] > ReadRequestQueue[MaxValue][9:0]) &&
                 !fsmWait[{ReadRequestQueue[i][40:39], ReadRequestQueue[i][38:37]}] &&
                 fsmIdle[{ReadRequestQueue[i][40:39], ReadRequestQueue[i][38:37]}]
                )begin
                    MaxValue = i[$clog2(CMDQUEUEDEPTH)-1:0];
                end else begin
                    MaxValue = MaxValue;
                end
            end
        end else begin
            for(int i = 0; i < WRITECMDQUEUEDEPTH; i++) begin
                if(!WriteReqQueFree[i] && (WriteRequestQueue[i][9:0] > WriteRequestQueue[MaxValue][9:0]) && 
                !fsmWait[{WriteRequestQueue[i][40:39], WriteRequestQueue[i][38:37]}] &&
                 fsmIdle[{WriteRequestQueue[i][40:39], WriteRequestQueue[i][38:37]}]
                )begin
                    MaxValue = i[$clog2(CMDQUEUEDEPTH)-1:0];
                end else begin
                    MaxValue = MaxValue;
                end
            end
        end
    end
    //  Checking Threshold in Aging, If THRESHOLD, PRIORITY chnaged to be 1   //
    always_comb begin 
        checkThreshold = 0;
        if(!WriteMode) begin
            // Read Request Serving
            for(int i = 0; i < READCMDQUEUEDEPTH; i++)begin
                if(!ReadReqQueFree[i] && (ReadRequestQueue[i][9:0] > THRESHOLD) &&
                !fsmWait[{ReadRequestQueue[i][40:39], ReadRequestQueue[i][38:37]}] &&
                 fsmIdle[{ReadRequestQueue[i][40:39], ReadRequestQueue[i][38:37]}]
                ) begin
                    checkThreshold = 1;
                end
            end
        end else begin
            // Write Request Serving
            for(int i= 0; i < WRITECMDQUEUEDEPTH; i++) begin
                if(!WriteReqQueFree[i] && (WriteRequestQueue[i][9:0] > THRESHOLD) &&
                !fsmWait[{WriteRequestQueue[i][40:39], WriteRequestQueue[i][38:37]}] &&
                 fsmIdle[{WriteRequestQueue[i][40:39], WriteRequestQueue[i][38:37]}]
                ) begin
                    checkThreshold = 1;
                end
            end
        end
    end

    //------------------------------------------------------------------------------
    //  FR-FCFS Final Selection
    //
    //  Priority Order:
    //      1) Requests beyond aging threshold
    //      2) Row-hit with short tCCD
    //      3) Row-hit with long tCCD
    //      4) Oldest request
    //
    //  - Determines final pop pointer.
    //  - Classifies PageHit / PageMiss / PageEmpty.
    //  - Decides auto-precharge behavior.
    //
    //------------------------------------------------------------------------------
    always_comb begin //FR-FCFS
        ReadPopPtr = 0;
        WritePopPtr = 0 ;
        checkAutoPrecharge  = 0;
        if(!WriteMode) begin 
            // Read Request Serving
            if(checkThreshold) begin                        // PRIORITY 1: Beyond Threshold, MOST AGING REQUEST
                ReadPopPtr = MaxValue;
                if(ReadOpenPagePolicyShort(MaxValue))begin
                    {PageHitT, PageMissT, PageEmptyT} =  4'b1000;
                end
                else if(ReadOpenPagePolicyLong(MaxValue)) begin
                    {PageHitT, PageMissT, PageEmptyT} = 4'b1100;
                end

                else if(OpenRowList[{ReadRequestQueue[MaxValue][40:39], ReadRequestQueue[MaxValue][38:37]}][15]) begin
                    {PageHitT, PageMissT, PageEmptyT} = 4'b0010;
                    checkAutoPrecharge = 1;                          // SPECULATIVE FOR MOST AGING REQUEST ON AUTO-PRECHARGE.
                                                                     // (TODO) Design Much More fancy scheme for eviction of entry in OpenPageList.
                end
                else begin
                    {PageHitT, PageMissT, PageEmptyT} = 4'b0001;
                end
            end
            else if(NextPageHitS) begin                     // PRIORITY 2: Case of PageHit & Short_tCCD
                ReadPopPtr = PageHitIndexS;
                {PageHitT, PageMissT, PageEmptyT} = 4'b1000;
            end
            else if(NextPageHitL) begin                     // PRIORITY 3: Case of PageHit & Long_tCCD
                ReadPopPtr = PageHitIndexL;
                {PageHitT, PageMissT, PageEmptyT} = 4'b1100;
            end
            else begin                                      // PRIORITY 4: Case of Aging-based Request Selection
                ReadPopPtr = MaxValue;
                if(OpenRowList[{ReadRequestQueue[MaxValue][40:39], ReadRequestQueue[MaxValue][38:37]}][15]) begin
                    {PageHitT, PageMissT, PageEmptyT}  =  4'b0010;
                end else begin
                    {PageHitT, PageMissT, PageEmptyT} =  4'b0001;
                end
            end
        end else begin
        // Write Request Serving
            if(checkThreshold) begin                        // PRIORITY 1: Beyond Threshold, MOST AGING REQUEST
                WritePopPtr = MaxValue;
                if(WriteOpenPagePolicyShort(MaxValue))begin
                    {PageHitT, PageMissT, PageEmptyT} =  4'b1000;
                end
                else if(WriteOpenPagePolicyLong(MaxValue)) begin
                    {PageHitT, PageMissT, PageEmptyT} = 4'b1100;
                end

                else if(OpenRowList[{WriteRequestQueue[MaxValue][40:39], WriteRequestQueue[MaxValue][38:37]}][15]) begin
                    {PageHitT, PageMissT, PageEmptyT} = 4'b0010;
                    checkAutoPrecharge = 1;
                end
                else begin
                    {PageHitT, PageMissT, PageEmptyT} = 4'b0001;
                end
            end
            else if(NextPageHitS) begin                     // PRIORITY 2: Case of PageHit & Short_tCCD
                WritePopPtr = PageHitIndexS;
                {PageHitT, PageMissT, PageEmptyT} = 4'b1000;
            end
            else if(NextPageHitL) begin                     // PRIORITY 3: Case of PageHit & Long_tCCD
                WritePopPtr = PageHitIndexL;
                {PageHitT, PageMissT, PageEmptyT} = 4'b1100;
            end
            else begin                                      // PRIORITY 4: Case of Aging-based Request Selection
                WritePopPtr = MaxValue;
                if(OpenRowList[{WriteRequestQueue[MaxValue][40:39], WriteRequestQueue[MaxValue][38:37]}][15]) begin
                    {PageHitT, PageMissT, PageEmptyT}  =  4'b0010;
                end else begin
                    {PageHitT, PageMissT, PageEmptyT} =  4'b0001;
                end
            end        
        end
    end
    
endmodule
